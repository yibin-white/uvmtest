`ifndef AXI_APB_SVH
`define AXI_APB_SVH


`include "axi_transfer.sv"
`include "apb_transfer.sv"
`include "axi_config.sv"

//master所有的头文件
`include "axi_driver.sv"
`include "apb_driver.sv"
`include "axi_sequencer.sv"
`include "axi_monitor.sv"

`include "axi_master_agent.sv"

`include "apb_monitor.sv"

`include "apb_slave_agent.sv"

//slave所有的头文件
`include "reference_model.sv"
`include "axi_scoreboard.sv"


//master头文件里面具体的实现方法



//env
`include "axi_env.sv" 

//sequence
`include "axi_apb_base_test_sequence.sv"       
`include "axi_sequence_addr.sv"
`include "axi_sequence_addr_burst.sv"
`include "axi_sequence_addr_read.sv"
`include "axi_sequence_addr_read_write.sv"
`include "virtual_sequence.sv"

`include "axi_addr_sequence_test.sv"
`include "axi_apb_base_test.sv"




   
`endif
